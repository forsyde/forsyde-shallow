library ieee;
use ieee.numeric_std.all;

package types is
  subtype int32 is signed(31 downto 0);  -- 32 bit integers 
end types;
